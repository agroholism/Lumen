﻿color-scheme='classic'
﻿color-scheme='oldstyle'